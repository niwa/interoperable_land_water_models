netcdf LUCI_output_netCDF_template {
dimensions:
	nrch = 532 ;
	time = UNLIMITED ; 
variables:
	int rchid(nrch) ;
		rchid:long_name = "identifier for stream reach" ;
	double time(time) ;
		time:standard_name = "time" ;
		time:units = "hours since 1970-01-01 0:00" ;
		time:axis = "T" ;
		time:calendar = "gregorian" ;
		time:bounds = "time_bnd" ;
		time:_FillValue = -9999. ;
	double ecotope_groundwater_recharge(time, nrch) ;
		ecotope_groundwater_recharge:description = "Groundwater recharge is baseflow plus interflow" ;
		ecotope_groundwater_recharge:standard_name = "(no standard name)" ;
		ecotope_groundwater_recharge:long_name = "Groundwater recharge (m3 s-1)" ;
		ecotope_groundwater_recharge:cdsm_name = "soil_water_sat-zone_top__recharge_volume_flux" ;
		ecotope_groundwater_recharge:units = "m3 s-1" ;
	double ecotope_fast_flow(time, nrch) ;
		ecotope_fast_flow:description = "The fast flow is throughflow plus overland flow" ;
		ecotope_fast_flow:standard_name = "(no standard name)" ;
		ecotope_fast_flow:cdsm_name = "land_surface_water__runoff_volume_flux" ;
		ecotope_fast_flow:long_name = "Fast flow (m3 s-1)" ;
		ecotope_fast_flow:units = "m3 s-1" ;
	double ecotope_gw_flow(time, nrch) ;
		ecotope_gw_flow:description = "The groundwater flow is baseflow plus interflow" ;
		ecotope_gw_flow:standard_name = "(no standard name)" ;
		ecotope_gw_flow:cdsm_name = "soil_water_unsat-zone__runoff_volume_flux" ;
		ecotope_gw_flow:long_name = "Groundwater flow (m3 s-1)" ;
		ecotope_gw_flow:units = "m3 s-1" ;

// global attributes:
		:title = "Output from rainfall runoff model" ;
		:institution = "Victoria University" ;
		:Conventions = "CF-1.7" ;
		:source = "LUCI" ;
		:comments = "Output from the Victoria University LUCI rainfall runoff model. The model outputs groundwater recharge and overland flow." ;
data:

 rchid = 15440662, 15440550, 15163382, 15440518, 15399270, 15440486, 
    15334790, 15440390, 15399094, 15440366, 15332702, 15440310, 15375494, 
    15440158, 15396294, 15439854, 15375350, 15439806, 15351446, 15439782, 
    15398374, 15439750, 15340126, 15439550, 15373990, 15439510, 15374166, 
    15439454, 15395262, 15439254, 15311390, 15439230, 15364846, 15438990, 
    15396038, 15438726, 15264086, 15438630, 15387430, 15438598, 15061126, 
    15438486, 15337846, 15438390, 15260262, 15438286, 15316342, 15438222, 
    15045574, 15307190, 15438102, 15318382, 15437982, 15425670, 15423798, 
    15437174, 15387125, 15375381, 15386709, 15361669, 15386573, 15347629, 
    15386141, 15316893, 15384685, 15373877, 15383685, 15292293, 15378493, 
    15383253, 15346805, 15367533, 15234821, 15313789, 15115133, 15375741, 
    15382469, 15374277, 15384125, 15275525, 15386389, 15386373, 15386965, 
    15330989, 15076525, 15082837, 15387357, 15354181, 15387453, 15074085, 
    15075205, 15388309, 15382317, 15388397, 15367661, 15388757, 15356005, 
    15388885, 15338205, 15389037, 15292021, 15396269, 15396093, 15399261, 
    15399109, 15399397, 15021813, 15020613, 15404453, 15404445, 15331422, 
    15315870, 15404501, 15377213, 15395822, 15307174, 15404509, 15370533, 
    15399102, 15396638, 15404517, 15274157, 15404525, 15376245, 15429958, 
    15430014, 15404405, 15395645, 15404597, 15394701, 15326300, 15302060, 
    15409453, 15336076, 15325716, 15197660, 15325628, 15317172, 15336084, 
    15249908, 15336100, 15165620, 15324796, 15315876, 15336108, 15283844, 
    15324212, 15316340, 15336124, 15282596, 15314212, 15336188, 15324196, 
    15283028, 15323412, 15374485, 15429902, 15424686, 15313596, 15323028, 
    15314180, 15291332, 15429854, 15396878, 15313636, 15207036, 15313572, 
    15274828, 15313500, 15247812, 15313292, 15210684, 15429694, 15372942, 
    15311708, 15312484, 15429550, 15336238, 15429502, 15423934, 15311916, 
    15312668, 15430318, 15363086, 15430518, 15334598, 15424654, 15430630, 
    15424470, 15423430, 15429030, 15366294, 15306772, 15307188, 15428726, 
    15374533, 15423894, 15348958, 15311052, 15307332, 15423726, 15423062, 
    15423526, 15423422, 15336228, 15295316, 15420446, 15419990, 15386093, 
    15421070, 15419270, 15419086, 15386029, 15314941, 15311668, 15274916, 
    15312052, 15133956, 15312908, 15336284, 15309484, 15282812, 15384133, 
    15310685, 15310372, 15272092, 15384005, 15377277, 15428486, 15394870, 
    15367213, 15375461, 15309060, 15285108, 15310388, 15292676, 15307468, 
    15302580, 15304484, 15296124, 15305460, 15308292, 15384741, 15338565, 
    15307732, 15308812, 15377653, 15361341, 15296476, 15303204, 15428126, 
    15319166, 15306556, 15258532, 15384165, 15338469, 15310204, 15322892, 
    15371965, 15427718, 15303428, 15250180, 15299972, 15301156, 15372869, 
    15365549, 15379957, 15343061, 15301916, 15282084, 15303548, 15249372, 
    15357085, 15357093, 15374749, 15369877, 15377325, 15311181, 15284268, 
    15218868, 15380613, 15357957, 15336292, 15287588, 15376117, 15329389, 
    15294580, 15255620, 15298692, 15293996, 15425606, 15425614, 15365645, 
    15333733, 15302108, 15263108, 15346101, 15344429, 15365973, 15354669, 
    15372117, 15354349, 15373957, 15372405, 15117124, 15189564, 15215044, 
    15359133, 15351301, 15301724, 15287836, 15311780, 15255588, 15364429, 
    15363893, 15356805, 15351813, 15129492, 15271268, 15369773, 15310461, 
    15297636, 15290308, 15304884, 15272372, 15311452, 15305324, 15367165, 
    15309181, 15374189, 15365557, 15365061, 15348837, 15302524, 15272036, 
    15359501, 15346997, 15363277, 15341165, 15365677, 15352013, 15365357, 
    15301525, 15290692, 15279996, 15361189, 15305061, 15287772, 15297668, 
    15395222, 15330374, 15300364, 15275284, 15362829, 15297341, 15287644, 
    15255972, 15354517, 15358413, 15342125, 15353093, 15289964, 15294020, 
    15425502, 15373214, 15388214, 15383622, 15284820, 15270708, 15356973, 
    15357909, 15359029, 15290149, 15361245, 15347445, 15360549, 15342445, 
    15357821, 15314525, 15363301, 15323373, 15297252, 15280932, 15395846, 
    15363006, 15359469, 15345885, 15288516, 15283620, 15361717, 15284989, 
    15346069, 15360637, 15394398, 15378582, 15361750, 15378966, 15357917, 
    15346701, 15279388, 15286500, 15290548, 15264652, 15425686, 15363262, 
    15379310, 15367942, 15352373, 15351821, 15430846, 15298198, 15355125, 
    15265781, 15292052, 15250236, 15349509, 15334765, 15383310, 15337606, 
    15347701, 15349045, 15366485, 15328109, 15436686, 15420278, 15310740, 
    15269844, 15302685, 15395869, 15424494, 15326390, 15354117, 15274277, 
    15290028, 15285708, 15365381, 15282709, 15338669, 15329197, 15339157, 
    15354613, 15338821, 15333309, 15350965, 15328893, 15384934, 15299078, 
    15421934, 15274862, 15276276, 15249844, 15136612, 15374150, 15353822, 
    15425846, 15344934, 15271068, 15264780, 15280516, 15260220, 15342245, 
    15335077, 15303076, 15268732, 15374374, 15315550, 15389438, 15372982, 
    15288940, 15275028, 15338381, 15314765, 15283364, 15234220, 15315109, 
    15308957, 15336885, 15320397, 15335869, 15268789, 15369190, 15285774, 
    15370830, 15361542, 15349053, 15306229, 15278924, 15256548, 15331421, 
    15315861, 15315077, 15325533, 15356702, 15326806, 15374110, 15295038, 
    15313989, 15324381, 15421286, 15305942, 15331669, 15311205, 15351445, 
    15292389, 15312086, 15296326, 15270532, 15222356, 15319789, 15307197, 
    15291612, 15243756, 15426086, 15321982, 15316525, 15277861, 15267188, 
    15301276, 15246196, 15252580, 15286292, 15306084, 15296877, 15297285, 
    15305021, 15248957, 15329158, 15319286, 15126053, 15249693, 15252981, 
    15130101 ;

 time = 1;
 }
